// adc_spi_frame_capture.v
//
// Generic framed SPI capture block.
//
// Goal (v1): provide a *usable* implementation with a stable interface for
// harness wiring + DV, without baking in ADS131M08-specific assumptions.
//
// Notes:
// - This block acts as a simple SPI master for read-only framed captures.
// - It generates SCLK + CS_N, drives MOSI low (NULL command).
// - It shifts in WORDS_PER_FRAME words of BITS_PER_WORD each from MISO.
// - Each captured word is right-justified into a 32-bit slot and packed into
//   frame_words_packed.
// - Packing convention: word 0 occupies bits [31:0], word 1 occupies [63:32], …
// - Bit order: MSB-first on the wire (first sampled bit becomes the MSB of the
//   word register).
//
// Timing model:
// - SCLK is generated by dividing clk with SCLK_DIV (must be >= 2).
// - CPOL/CPHA are parameterized; default matches ADS131M08 mode (CPOL=0, CPHA=1)
//   per project spec.
//
`default_nettype none

module adc_spi_frame_capture #(
    parameter int unsigned BITS_PER_WORD   = 24,
    parameter int unsigned WORDS_PER_FRAME = 9,

    // Divide ratio for SCLK relative to clk. SCLK toggles every SCLK_DIV cycles.
    // => full SCLK period = 2*SCLK_DIV cycles.
    parameter int unsigned SCLK_DIV        = 4,

    // SPI mode select
    parameter bit          CPOL            = 1'b0,
    parameter bit          CPHA            = 1'b1
) (
    input  wire                          clk,
    input  wire                          rst,

    // Start capture for one frame (pulse)
    input  wire                          start,

    // SPI pins (direction is from our SoC perspective)
    output wire                          adc_sclk,
    output wire                          adc_cs_n,
    output wire                          adc_mosi,
    input  wire                          adc_miso,

    // Frame result
    output wire                          frame_valid,
    output wire [32*WORDS_PER_FRAME-1:0]  frame_words_packed,

    output wire                          busy
);

    // -------------------------
    // Parameter sanity
    // -------------------------
    initial begin
        if (BITS_PER_WORD == 0) begin
            $error("adc_spi_frame_capture: BITS_PER_WORD must be > 0");
        end
        if (WORDS_PER_FRAME == 0) begin
            $error("adc_spi_frame_capture: WORDS_PER_FRAME must be > 0");
        end
        if (BITS_PER_WORD > 32) begin
            $error("adc_spi_frame_capture: BITS_PER_WORD must be <= 32 for 32b packing");
        end
        if (SCLK_DIV < 2) begin
            $error("adc_spi_frame_capture: SCLK_DIV must be >= 2");
        end
    end

    // -------------------------
    // Internal regs
    // -------------------------
    localparam int unsigned WORD_BITS_W = (BITS_PER_WORD < 2) ? 1 : $clog2(BITS_PER_WORD);
    localparam int unsigned WORDS_W     = (WORDS_PER_FRAME < 2) ? 1 : $clog2(WORDS_PER_FRAME);

    reg                         busy_r;
    reg                         frame_valid_r;

    reg                         cs_n_r;
    reg                         sclk_r;
    reg [$clog2(SCLK_DIV)-1:0]   div_ctr_r;

    reg [WORD_BITS_W:0]          bit_idx_r;   // 0..BITS_PER_WORD
    reg [WORDS_W:0]              word_idx_r;  // 0..WORDS_PER_FRAME
    reg [BITS_PER_WORD-1:0]      word_shift_r;
    reg [32*WORDS_PER_FRAME-1:0] frame_words_r;

    // Track whether the upcoming toggle is a leading edge (low->high) or trailing.
    wire next_sclk = ~sclk_r;
    wire is_leading_edge  = (sclk_r == 1'b0) && (next_sclk == 1'b1);
    wire is_trailing_edge = (sclk_r == 1'b1) && (next_sclk == 1'b0);

    // For CPOL=1, the notion of leading/trailing relative to idle flips.
    // Define "leading" as the first edge away from idle, and "trailing" as return-to-idle.
    wire sclk_idle = CPOL;
    wire leaving_idle  = (sclk_r == sclk_idle) && (next_sclk != sclk_idle);
    wire returning_idle = (sclk_r != sclk_idle) && (next_sclk == sclk_idle);

    wire is_spi_leading  = leaving_idle;
    wire is_spi_trailing = returning_idle;

    // Sample edge selection:
    // CPHA=0 => sample on leading edge
    // CPHA=1 => sample on trailing edge
    wire sample_on_toggle = (CPHA == 1'b0) ? is_spi_leading : is_spi_trailing;

    // -------------------------
    // Outputs
    // -------------------------
    assign adc_cs_n          = cs_n_r;
    assign adc_sclk          = sclk_r;
    assign adc_mosi          = 1'b0;  // NULL command in v1

    assign frame_valid       = frame_valid_r;
    assign frame_words_packed = frame_words_r;
    assign busy              = busy_r;

    // -------------------------
    // Capture FSM (single-state busy/idle)
    // -------------------------
    always @(posedge clk) begin
        if (rst) begin
            busy_r        <= 1'b0;
            frame_valid_r <= 1'b0;
            cs_n_r        <= 1'b1;
            sclk_r        <= sclk_idle;
            div_ctr_r     <= '0;

            bit_idx_r     <= '0;
            word_idx_r    <= '0;
            word_shift_r  <= '0;
            frame_words_r <= '0;
        end else begin
            frame_valid_r <= 1'b0; // default: pulse

            if (!busy_r) begin
                cs_n_r    <= 1'b1;
                sclk_r    <= sclk_idle;
                div_ctr_r <= '0;

                bit_idx_r  <= '0;
                word_idx_r <= '0;
                word_shift_r <= '0;

                if (start) begin
                    busy_r        <= 1'b1;
                    cs_n_r        <= 1'b0;
                    // Clear output container at start-of-frame.
                    frame_words_r <= '0;
                end
            end else begin
                // busy_r == 1
                // Generate SCLK toggles with divider.
                if (div_ctr_r == SCLK_DIV-1) begin
                    div_ctr_r <= '0;
                    sclk_r    <= next_sclk;

                    if (sample_on_toggle) begin
                        // Shift MSB-first: first sampled bit becomes MSB of word.
                        word_shift_r <= {word_shift_r[BITS_PER_WORD-2:0], adc_miso};
                        bit_idx_r    <= bit_idx_r + 1'b1;

                        if (bit_idx_r == BITS_PER_WORD-1) begin
                            // Completed a word.
                            // Right-justify into 32b slot (zero-extend).
                            frame_words_r[32*word_idx_r +: 32] <= {{(32-BITS_PER_WORD){1'b0}}, {word_shift_r[BITS_PER_WORD-2:0], adc_miso}};

                            bit_idx_r    <= '0;
                            word_shift_r <= '0;
                            word_idx_r   <= word_idx_r + 1'b1;

                            if (word_idx_r == WORDS_PER_FRAME-1) begin
                                // Completed the last word; end capture.
                                busy_r        <= 1'b0;
                                cs_n_r        <= 1'b1;
                                sclk_r        <= sclk_idle;
                                frame_valid_r <= 1'b1;
                            end
                        end
                    end
                end else begin
                    div_ctr_r <= div_ctr_r + 1'b1;
                end
            end
        end
    end

endmodule

`default_nettype wire
